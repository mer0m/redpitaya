library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

Entity wb_nco_counter is 
    generic(
		COUNTER_SIZE : natural := 32;
        id        : natural := 1;
        wb_size   : natural := 16 -- Data port size for wishbone
    );
    port 
    (
		-- Syscon signals
		reset     : in std_logic ;
		clk       : in std_logic ;
		-- Wishbone signals
		wbs_add       : in std_logic_vector(1 downto 0);
		wbs_write     : in std_logic ;
		wbs_writedata : in std_logic_vector( wb_size-1 downto 0);
		wbs_read     : in std_logic ;
		wbs_readdata  : out std_logic_vector( wb_size-1 downto 0);
		pinc_sw_o 		: out std_logic;
		poff_sw_o 		: out std_logic;
		cpt_off_o	: out std_logic_vector(COUNTER_SIZE-1 downto 0);
		cpt_step_o : out std_logic_vector(COUNTER_SIZE-1 downto 0)
    );
end entity wb_nco_counter;


-----------------------------------------------------------------------
Architecture wb_nco_counter_1 of wb_nco_counter is
-----------------------------------------------------------------------
	constant REG_ID     : std_logic_vector := "00";
	constant REG_PINC 	: std_logic_vector :="01";
	constant REG_POFF 	: std_logic_vector :="10";
	constant REG_CTRL 	: std_logic_vector :="11";
	signal cpt_step_s 	: std_logic_vector(31 downto 0);
	signal cpt_off_s 	: std_logic_vector(31 downto 0);
	signal poff_sw_s	: std_logic;
	signal pinc_sw_s	: std_logic;
	signal readdata_s 	: std_logic_vector(wb_size-1 downto 0);
begin
	wbs_readdata <= readdata_s;
	cpt_step_o <= cpt_step_s(COUNTER_SIZE-1 downto 0);
	cpt_off_o <= cpt_off_s(COUNTER_SIZE-1 downto 0);
	pinc_sw_o <= pinc_sw_s;
	poff_sw_o <= poff_sw_s;
	-- manage register
	write_bloc : process(clk, reset)   -- write DEPUIS l'iMx
	begin
		 if reset = '1' then 
			cpt_step_s <= x"0A3D70A3";--(COUNTER_SIZE-1 downto 5 => '0')&"11000";--(others =>'0' );
			cpt_off_s <= (others => '0');
			pinc_sw_s <= '1';
			poff_sw_s <= '1';
		 elsif rising_edge(clk) then
			cpt_step_s <= cpt_step_s;
			cpt_off_s <= cpt_off_s;
			pinc_sw_s <= pinc_sw_s;
			poff_sw_s <= poff_sw_s;
			if (wbs_write = '1' ) then
				case wbs_add is
				when REG_PINC =>
					cpt_step_s <= wbs_writedata;
				when REG_POFF =>
					cpt_off_s <= wbs_writedata;
				when REG_CTRL =>
					pinc_sw_s <= wbs_writedata(0);
					poff_sw_s <= wbs_writedata(1);
				when others =>
				end case;
			  end if;
		 end if;
	end process write_bloc;

	read_bloc : process(clk, reset)
	begin
		if reset = '1' then
			readdata_s <= (others => '0');
		elsif rising_edge(clk) then
			readdata_s <= readdata_s;
			if (wbs_read = '1') then
				case wbs_add is
				when REG_ID =>
					 readdata_s <= std_logic_vector(to_unsigned(id,wb_size));
				when REG_PINC =>
					readdata_s <= cpt_step_s;
				when REG_POFF =>
					readdata_s <= cpt_off_s;
				when REG_CTRL =>
					readdata_s <= (wb_size-1 downto 2 => '0')&poff_sw_s&pinc_sw_s;
				when others =>
					readdata_s <= (others => '0');
				end case;
			end if;
		end if;
	end process read_bloc;

end architecture wb_nco_counter_1;

